module InstructionMemory(PC, InstructOut);
	input[31:0] PC;
	reg [31:0] Instruction[31:0];
	output [31:0] InstructOut;
	always@(PC) begin
		if(PC == 32'b00000000000000000000000000000000) begin
			/*//R[0]!
			Instruction[0] = 32'b010011_00000_000000000000000000000;  //R[0] = In
			Instruction[1] = 32'b010100_00000_000000000000000000000; //Out[R[0]]
 			Instruction[2] = 32'b000110_00001_000000000000000000001;  //R[1] = 1
			Instruction[3] = 32'b000110_01000_000000000000000000101;  //R[8] = 5
			Instruction[4] = 32'b000100_00001_00010_0000000000000000; //R[2] = R[1]
			//R[3] = R[1] * R[2]
			Instruction[5] = 32'b000100_00001_00110_0000000000000000; //R[6] = R[1]
			Instruction[6] = 32'b000110_01001_000000000000000000000;  //R[9] = 0
			Instruction[7] = 32'b000110_00100_000000000000000000001;  //R[4] = 1
			Instruction[8] = 32'b000110_00101_000000000000000001010;  //R[5] = 10 -> posição da da soma
			Instruction[9] = 32'b000110_00011_000000000000000000000;  //R[3] = 0
			//multiplicacao
			Instruction[10]= 32'b000001_00011_00010_00011_00000000000;//R[3] = R[2] + R[3]
			Instruction[11]= 32'b000010_00110_00100_00110_00000000000;//R[6] = R[6] - R[4]
			Instruction[12]= 32'b001111_00110_01001_00101_00000000000;//Se R[6] > R[9] -> PC = R[5] senão PC = PC++
			//condicional
			Instruction[13]= 32'b000100_00011_00010_0000000000000000; //R[2] = R[3]
			Instruction[14]= 32'b010100_00010_000000000000000000000; //Out[R[2]]
			Instruction[15]= 32'b000001_00001_00100_00001_00000000000;//R[1] = R[4] +R[1]
			Instruction[16]= 32'b001111_00000_00001_01000_00000000000;//Se R[0] > R[1] -> PC = R[8] senão PC = PC++
			Instruction[17]= 32'b000000_00000000000000000000000000; //NOP
			Instruction[18]= 32'b001101_00000_00001_01000_00000000000;//Se R[0] == R[1] -> PC = R[8] senão PC = PC++
			Instruction[19]= 32'b000101_00101_00010_0000000000000000; //Mem[R[5]] = R[2]
			Instruction[20]= 32'b000000_00000000000000000000000000; //NOP
			Instruction[21]= 32'b000011_00101_01111_0000000000000000;//R[15] = Mem[R[5]]
			Instruction[22]= 32'b010100_01111_000000000000000000000; //Out[R[15]]
			Instruction[23]= 32'b111111_00000000000000000000000000; //halt
			*/
			
			/*
			//Algoritmo teste
			
			Instruction[0] = 32'b000110_00000_000000000000000000001;			//R[0] = 1
			Instruction[1] = 32'b001100_00000_00000_00001_00001_000000; 	//R[1] = R[0] << 1 = 2
			Instruction[2] = 32'b001011_00001_00000_00010_00001_000000;		//R[2] = R[1] >> 1 = 1
			Instruction[3] = 32'b000001_00001_00010_00100_00000000000;		//R[4] = R[2] + R[1] = 3
			Instruction[4] = 32'b000010_00001_00010_00011_00000000000;     //R[3] = R[1] - R[2] = 1
			Instruction[5] = 32'b001101_00011_00100_00100_00000000000;		//Se R[3] == R[4] -> PC = R[4] senao PC++
			Instruction[6] = 32'b000110_00101_000000000000000000111;			//R[5] = 7
			Instruction[7] = 32'b000001_00000_00010_00000_00000000000;		//R[0] = R[2] + R[0]
			Instruction[8] = 32'b001110_00000_00100_00101_00000000000;		//Se R[0] != R[4] -> PC = R[5] senao PC++
			Instruction[9] = 32'b001000_00000_00000_0000_000000000000;		//R[0] = R[0] | R[0]
			Instruction[10]= 32'b001001_00000_00000_0000000000000000;		//R[0] = ~R[0]
			Instruction[11]= 32'b000111_00000_00000_00000_00000000000;		//R[0] = R[0] & R[0]
			Instruction[12]= 32'b010001_0000000000_00000_00000001110;		//jump 14
			Instruction[13]= 32'b111111_00000000000000000000000000;			//halt
			Instruction[14]= 32'b001010_00000_00000_00001_00000000000;		//R[0] = R[0] xor R[0]
			Instruction[15]= 32'b010100_00000_000000000000000000000; 		//Out[R[0]]
			Instruction[16]= 32'b010010_00001_000000000000000000000;			//Jr R[1]
			*/
			
			//Teste Instrucoes
			
			Instruction[0] = 32'b000110_00000_000000000000000000001;			// li R[0] 1
			Instruction[1] = 32'b000110_00001_000000000000000000011;			// li R[1] 3
			Instruction[2] = 32'b000000_00000000000000000000000000;			// nop
			Instruction[3] = 32'b000001_00000_00001_00010_0000000000;		// add R[0] R[1] R[2]
			Instruction[4] = 32'b000010_00000_00001_00010_0000000000;		// sub R[0] R[1] R[2]
			Instruction[5] = 32'b000011_00000_00001_000000000000000;			// lw R[0] R[1]
			Instruction[6] = 32'b000100_00010_00100_000000000000000;			// mov R[2] R[4]
			Instruction[7] = 32'b000101_00000_00101_000000000000000;			// sw R[0] R[5]
			Instruction[8] = 32'b000110_00110_00000000000000000000;			// li R[6] 0
			Instruction[9] = 32'b000111_00000_00110_00111_0000000000;		// and R[0] R[6] R[7]
			Instruction[10]= 32'b001000_00000_00110_00111_0000000000;		// or R[0] R[6] R[7]
			Instruction[11]= 32'b001001_00000_00111_000000000000000;			// not R[0] R[7]
			Instruction[12]= 32'b001010_00111_00111_00111_0000000000;		// xor R[7] R[7] R[7]
			Instruction[13]= 32'b001011_00001_00000_00111_00001_00000;		// sll R[1] R[7] 1
			Instruction[14]= 32'b001100_00001_00000_00111_00001_00000;		// srl R[1] R[7] 1
			Instruction[15]= 32'b000110_00111_000000000000000000001;			// li R[7] 1
			Instruction[16]= 32'b000110_01000_000000000000000000010;			// li R[8] 2
			Instruction[17]= 32'b001101_00000_00000_00000_00000000000;		// 
			Instruction[]= 32'b001101
			
			
		end
	end
	assign InstructOut = Instruction[PC];
endmodule

